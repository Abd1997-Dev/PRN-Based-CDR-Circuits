`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 20.04.2023 10:11:29
// Design Name: 
// Module Name: D_ff
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module D_ff(input d, clk, rst, output reg q);
 always @ (posedge clk) begin
 if (rst) q <= 0;
 else q <= d;
 end
endmodule


/*module d_ff(input din, clk, rst, output reg dout);
 always @ (posedge clk) begin
 if (rst) dout <= 0;
 else dout <= din;
 end
endmodule*/
